// Parameters used to define the data format and locations of fields within the ethernet header




